//CALIPTRA fuse data is in a memory space mapped from address 0x100 as an example
`define CALIPTRA_UDS_SEED_0                            32'h0000100
`define CALIPTRA_UDS_SEED_0_MASK                       32'hffffffff
`define CALIPTRA_UDS_SEED_1                            32'h0000104
`define CALIPTRA_UDS_SEED_1_MASK                       32'hffffffff
`define CALIPTRA_UDS_SEED_2                            32'h0000108
`define CALIPTRA_UDS_SEED_2_MASK                       32'hffffffff
`define CALIPTRA_UDS_SEED_3                            32'h000010C
`define CALIPTRA_UDS_SEED_3_MASK                       32'hffffffff
`define CALIPTRA_UDS_SEED_4                            32'h0000110
`define CALIPTRA_UDS_SEED_4_MASK                       32'hffffffff
`define CALIPTRA_UDS_SEED_5                            32'h0000114
`define CALIPTRA_UDS_SEED_5_MASK                       32'hffffffff
`define CALIPTRA_UDS_SEED_6                            32'h0000118
`define CALIPTRA_UDS_SEED_6_MASK                       32'hffffffff
`define CALIPTRA_UDS_SEED_7                            32'h000011c
`define CALIPTRA_UDS_SEED_7_MASK                       32'hffffffff
`define CALIPTRA_UDS_SEED_8                            32'h0000120
`define CALIPTRA_UDS_SEED_8_MASK                       32'hffffffff
`define CALIPTRA_UDS_SEED_9                            32'h0000124
`define CALIPTRA_UDS_SEED_9_MASK                       32'hffffffff
`define CALIPTRA_UDS_SEED_10                           32'h0000128
`define CALIPTRA_UDS_SEED_10_MASK                      32'hffffffff
`define CALIPTRA_UDS_SEED_11                           32'h000012c
`define CALIPTRA_UDS_SEED_11_MASK                      32'hffffffff
`define CALIPTRA_FIELD_ENTROPY_0                       32'h0000130
`define CALIPTRA_FIELD_ENTROPY_0_MASK                  32'hffffffff
`define CALIPTRA_FIELD_ENTROPY_1                       32'h0000134
`define CALIPTRA_FIELD_ENTROPY_1_MASK                  32'hffffffff
`define CALIPTRA_FIELD_ENTROPY_2                       32'h0000138
`define CALIPTRA_FIELD_ENTROPY_2_MASK                  32'hffffffff
`define CALIPTRA_FIELD_ENTROPY_3                       32'h000013c
`define CALIPTRA_FIELD_ENTROPY_3_MASK                  32'hffffffff
`define CALIPTRA_FIELD_ENTROPY_4                       32'h0000140
`define CALIPTRA_FIELD_ENTROPY_4_MASK                  32'hffffffff
`define CALIPTRA_FIELD_ENTROPY_5                       32'h0000144
`define CALIPTRA_FIELD_ENTROPY_5_MASK                  32'hffffffff
`define CALIPTRA_FIELD_ENTROPY_6                       32'h0000148
`define CALIPTRA_FIELD_ENTROPY_6_MASK                  32'hffffffff
`define CALIPTRA_FIELD_ENTROPY_7                       32'h000014c
`define CALIPTRA_FIELD_ENTROPY_7_MASK                  32'hffffffff
`define CALIPTRA_KEY_MANIFEST_PK_HASH_0                32'h0000150
`define CALIPTRA_KEY_MANIFEST_PK_HASH_0_MASK           32'hffffffff
`define CALIPTRA_KEY_MANIFEST_PK_HASH_1                32'h0000154
`define CALIPTRA_KEY_MANIFEST_PK_HASH_1_MASK           32'hffffffff
`define CALIPTRA_KEY_MANIFEST_PK_HASH_2                32'h0000158
`define CALIPTRA_KEY_MANIFEST_PK_HASH_2_MASK           32'hffffffff
`define CALIPTRA_KEY_MANIFEST_PK_HASH_3                32'h000015c
`define CALIPTRA_KEY_MANIFEST_PK_HASH_3_MASK           32'hffffffff
`define CALIPTRA_KEY_MANIFEST_PK_HASH_4                32'h0000160
`define CALIPTRA_KEY_MANIFEST_PK_HASH_4_MASK           32'hffffffff
`define CALIPTRA_KEY_MANIFEST_PK_HASH_5                32'h0000164
`define CALIPTRA_KEY_MANIFEST_PK_HASH_5_MASK           32'hffffffff
`define CALIPTRA_KEY_MANIFEST_PK_HASH_6                32'h0000168
`define CALIPTRA_KEY_MANIFEST_PK_HASH_6_MASK           32'hffffffff
`define CALIPTRA_KEY_MANIFEST_PK_HASH_7                32'h000016c
`define CALIPTRA_KEY_MANIFEST_PK_HASH_7_MASK           32'hffffffff
`define CALIPTRA_KEY_MANIFEST_PK_HASH_8                32'h0000170
`define CALIPTRA_KEY_MANIFEST_PK_HASH_8_MASK           32'hffffffff
`define CALIPTRA_KEY_MANIFEST_PK_HASH_9                32'h0000174
`define CALIPTRA_KEY_MANIFEST_PK_HASH_9_MASK           32'hffffffff
`define CALIPTRA_KEY_MANIFEST_PK_HASH_10               32'h0000178
`define CALIPTRA_KEY_MANIFEST_PK_HASH_10_MASK          32'hffffffff
`define CALIPTRA_KEY_MANIFEST_PK_HASH_11               32'h000017c
`define CALIPTRA_KEY_MANIFEST_PK_HASH_11_MASK          32'hffffffff
`define CALIPTRA_OWNER_PK_HASH_0                       32'h0000180
`define CALIPTRA_OWNER_PK_HASH_0_MASK                  32'hffffffff
`define CALIPTRA_OWNER_PK_HASH_1                       32'h0000184
`define CALIPTRA_OWNER_PK_HASH_1_MASK                  32'hffffffff
`define CALIPTRA_OWNER_PK_HASH_2                       32'h0000188
`define CALIPTRA_OWNER_PK_HASH_2_MASK                  32'hffffffff
`define CALIPTRA_OWNER_PK_HASH_3                       32'h000018c
`define CALIPTRA_OWNER_PK_HASH_3_MASK                  32'hffffffff
`define CALIPTRA_OWNER_PK_HASH_4                       32'h0000190
`define CALIPTRA_OWNER_PK_HASH_4_MASK                  32'hffffffff
`define CALIPTRA_OWNER_PK_HASH_5                       32'h0000194
`define CALIPTRA_OWNER_PK_HASH_5_MASK                  32'hffffffff
`define CALIPTRA_OWNER_PK_HASH_6                       32'h0000198
`define CALIPTRA_OWNER_PK_HASH_6_MASK                  32'hffffffff
`define CALIPTRA_OWNER_PK_HASH_7                       32'h000019c
`define CALIPTRA_OWNER_PK_HASH_7_MASK                  32'hffffffff
`define CALIPTRA_OWNER_PK_HASH_8                       32'h00001a0
`define CALIPTRA_OWNER_PK_HASH_8_MASK                  32'hffffffff
`define CALIPTRA_OWNER_PK_HASH_9                       32'h00001a4
`define CALIPTRA_OWNER_PK_HASH_9_MASK                  32'hffffffff
`define CALIPTRA_OWNER_PK_HASH_10                      32'h00001a8
`define CALIPTRA_OWNER_PK_HASH_10_MASK                 32'hffffffff
`define CALIPTRA_OWNER_PK_HASH_11                      32'h00001ac
`define CALIPTRA_OWNER_PK_HASH_11_MASK                 32'hffffffff
`define CALIPTRA_KEY_MANIFEST_SVN                      32'h00001b0
`define CALIPTRA_KEY_MANIFEST_SVN_MASK                 32'hffffffff
`define CALIPTRA_RUNTIME_SVN_0                         32'h00001b4
`define CALIPTRA_RUNTIME_SVN_0_MASK                    32'hffffffff
`define CALIPTRA_RUNTIME_SVN_1                         32'h00001b8
`define CALIPTRA_RUNTIME_SVN_1_MASK                    32'hffffffff
`define CALIPTRA_RUNTIME_SVN_2                         32'h00001bc
`define CALIPTRA_RUNTIME_SVN_2_MASK                    32'hffffffff
`define CALIPTRA_RUNTIME_SVN_3                         32'h00001c0
`define CALIPTRA_RUNTIME_SVN_3_MASK                    32'hffffffff
`define CALIPTRA_PUBLIC_SERIAL_NUMBER_0                32'h00001c4
`define CALIPTRA_PUBLIC_SERIAL_NUMBER_0_MASK           32'hffffffff
`define CALIPTRA_PUBLIC_SERIAL_NUMBER_1                32'h00001c8
`define CALIPTRA_PUBLIC_SERIAL_NUMBER_1_MASK           32'hffffffff
`define CALIPTRA_PUBLIC_SERIAL_NUMBER_2                32'h00001cc
`define CALIPTRA_PUBLIC_SERIAL_NUMBER_2_MASK           32'hffffffff
`define CALIPTRA_PUBLIC_SERIAL_NUMBER_3                32'h00001d0
`define CALIPTRA_PUBLIC_SERIAL_NUMBER_3_MASK           32'hffffffff
`define CALIPTRA_LMS_KEY_REVOKE_MASK                   32'h00001d4
`define CALIPTRA_LMS_KEY_REVOKE_MASK_MASK              32'hffffffff
`define CALIPTRA_FPF_TRNG_0                            32'h00001d8
`define CALIPTRA_FPF_TRNG_0_MASK                       32'hffffffff
`define CALIPTRA_FPF_TRNG_1                            32'h00001dc
`define CALIPTRA_FPF_TRNG_1_MASK                       32'h0000ffff
`define CALIPTRA_FPF_WDT                               32'h00001dc
`define CALIPTRA_FPF_WDT_MASK                          32'h00030000
`define CALIPTRA_HW_ID                                 32'h00001dc
`define CALIPTRA_HW_ID_MASK                            32'h03FC0000
`define CALIPTRA_ANTI_ROLLBACK_DISABLE                 32'h00001e0
`define CALIPTRA_ANTI_ROLLBACK_DISABLE_MASK            32'h00000001
`define CALIPTRA_KEY_MANIFEST_PK_HASH_MASK             32'h00001e0
`define CALIPTRA_KEY_MANIFEST_PK_HASH_MASK_MASK        32'h0000001E
`define CALIPTRA_LMS_VERIFY_ENABLE                     32'h00001e0
`define CALIPTRA_LMS_VERIFY_ENABLE_MASK                32'h00000020
`define CALIPTRA_IDEVID_CSR_REQUEST                    32'h00001e0
`define CALIPTRA_IDEVID_CSR_REQUEST_MASK               32'h00000040
`define CALIPTRA_CERT_ATTRIB_RATS                      32'h00001e0
`define CALIPTRA_CERT_ATTRIB_RATS_MASK                 32'h00000080
`define CALIPTRA_SET_FUSE_DONE                         32'h00001e0
`define CALIPTRA_SET_FUSE_DONE_MASK                    32'h00000100
