module caliptra_fdm_lut_fetch
  import fuse_lut_pkg::*;
(
  input                                  i_clk,
  input                                  i_readen,
  input  [$clog2(LUT_ENTRIES)-1:0]       i_raddr,
  output [$bits(fuse_lut_element_t)-1:0] o_rdata
);
  
  parameter fuse_lut_element_t FUSE_LUT[LUT_ENTRIES] = '{
    {`CALIPTRA_UDS_SEED_0_MASK,                 `CALIPTRA_UDS_SEED_0,                 `CLP_SOC_IFC_REG_FUSE_UDS_SEED_0},
    {`CALIPTRA_UDS_SEED_1_MASK,                 `CALIPTRA_UDS_SEED_1,                 `CLP_SOC_IFC_REG_FUSE_UDS_SEED_1},
    {`CALIPTRA_UDS_SEED_2_MASK,                 `CALIPTRA_UDS_SEED_2,                 `CLP_SOC_IFC_REG_FUSE_UDS_SEED_2},
    {`CALIPTRA_UDS_SEED_3_MASK,                 `CALIPTRA_UDS_SEED_3,                 `CLP_SOC_IFC_REG_FUSE_UDS_SEED_3},
    {`CALIPTRA_UDS_SEED_4_MASK,                 `CALIPTRA_UDS_SEED_4,                 `CLP_SOC_IFC_REG_FUSE_UDS_SEED_4},
    {`CALIPTRA_UDS_SEED_5_MASK,                 `CALIPTRA_UDS_SEED_5,                 `CLP_SOC_IFC_REG_FUSE_UDS_SEED_5},
    {`CALIPTRA_UDS_SEED_6_MASK,                 `CALIPTRA_UDS_SEED_6,                 `CLP_SOC_IFC_REG_FUSE_UDS_SEED_6},
    {`CALIPTRA_UDS_SEED_7_MASK,                 `CALIPTRA_UDS_SEED_7,                 `CLP_SOC_IFC_REG_FUSE_UDS_SEED_7},
    {`CALIPTRA_UDS_SEED_8_MASK,                 `CALIPTRA_UDS_SEED_8,                 `CLP_SOC_IFC_REG_FUSE_UDS_SEED_8},
    {`CALIPTRA_UDS_SEED_9_MASK,                 `CALIPTRA_UDS_SEED_9,                 `CLP_SOC_IFC_REG_FUSE_UDS_SEED_9},
    {`CALIPTRA_UDS_SEED_10_MASK,                `CALIPTRA_UDS_SEED_10,                `CLP_SOC_IFC_REG_FUSE_UDS_SEED_10},
    {`CALIPTRA_UDS_SEED_11_MASK,                `CALIPTRA_UDS_SEED_11,                `CLP_SOC_IFC_REG_FUSE_UDS_SEED_11},
    {`CALIPTRA_FIELD_ENTROPY_0_MASK,            `CALIPTRA_FIELD_ENTROPY_0,            `CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_0},
    {`CALIPTRA_FIELD_ENTROPY_1_MASK,            `CALIPTRA_FIELD_ENTROPY_1,            `CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_1},
    {`CALIPTRA_FIELD_ENTROPY_2_MASK,            `CALIPTRA_FIELD_ENTROPY_2,            `CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_2},
    {`CALIPTRA_FIELD_ENTROPY_3_MASK,            `CALIPTRA_FIELD_ENTROPY_3,            `CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_3},
    {`CALIPTRA_FIELD_ENTROPY_4_MASK,            `CALIPTRA_FIELD_ENTROPY_4,            `CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_4},
    {`CALIPTRA_FIELD_ENTROPY_5_MASK,            `CALIPTRA_FIELD_ENTROPY_5,            `CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_5},
    {`CALIPTRA_FIELD_ENTROPY_6_MASK,            `CALIPTRA_FIELD_ENTROPY_6,            `CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_6},
    {`CALIPTRA_FIELD_ENTROPY_7_MASK,            `CALIPTRA_FIELD_ENTROPY_7,            `CLP_SOC_IFC_REG_FUSE_FIELD_ENTROPY_7},
    {`CALIPTRA_KEY_MANIFEST_PK_HASH_0_MASK,     `CALIPTRA_KEY_MANIFEST_PK_HASH_0,     `CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_0},
    {`CALIPTRA_KEY_MANIFEST_PK_HASH_1_MASK,     `CALIPTRA_KEY_MANIFEST_PK_HASH_1,     `CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_1},
    {`CALIPTRA_KEY_MANIFEST_PK_HASH_2_MASK,     `CALIPTRA_KEY_MANIFEST_PK_HASH_2,     `CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_2},
    {`CALIPTRA_KEY_MANIFEST_PK_HASH_3_MASK,     `CALIPTRA_KEY_MANIFEST_PK_HASH_3,     `CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_3},
    {`CALIPTRA_KEY_MANIFEST_PK_HASH_4_MASK,     `CALIPTRA_KEY_MANIFEST_PK_HASH_4,     `CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_4},
    {`CALIPTRA_KEY_MANIFEST_PK_HASH_5_MASK,     `CALIPTRA_KEY_MANIFEST_PK_HASH_5,     `CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_5},
    {`CALIPTRA_KEY_MANIFEST_PK_HASH_6_MASK,     `CALIPTRA_KEY_MANIFEST_PK_HASH_6,     `CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_6},
    {`CALIPTRA_KEY_MANIFEST_PK_HASH_7_MASK,     `CALIPTRA_KEY_MANIFEST_PK_HASH_7,     `CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_7},
    {`CALIPTRA_KEY_MANIFEST_PK_HASH_8_MASK,     `CALIPTRA_KEY_MANIFEST_PK_HASH_8,     `CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_8},
    {`CALIPTRA_KEY_MANIFEST_PK_HASH_9_MASK,     `CALIPTRA_KEY_MANIFEST_PK_HASH_9,     `CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_9},
    {`CALIPTRA_KEY_MANIFEST_PK_HASH_10_MASK,    `CALIPTRA_KEY_MANIFEST_PK_HASH_10,    `CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_10},
    {`CALIPTRA_KEY_MANIFEST_PK_HASH_11_MASK,    `CALIPTRA_KEY_MANIFEST_PK_HASH_11,    `CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_11},
    {`CALIPTRA_OWNER_PK_HASH_0_MASK,            `CALIPTRA_OWNER_PK_HASH_0,            `CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_0},
    {`CALIPTRA_OWNER_PK_HASH_1_MASK,            `CALIPTRA_OWNER_PK_HASH_1,            `CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_1},
    {`CALIPTRA_OWNER_PK_HASH_2_MASK,            `CALIPTRA_OWNER_PK_HASH_2,            `CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_2},
    {`CALIPTRA_OWNER_PK_HASH_3_MASK,            `CALIPTRA_OWNER_PK_HASH_3,            `CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_3},
    {`CALIPTRA_OWNER_PK_HASH_4_MASK,            `CALIPTRA_OWNER_PK_HASH_4,            `CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_4},
    {`CALIPTRA_OWNER_PK_HASH_5_MASK,            `CALIPTRA_OWNER_PK_HASH_5,            `CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_5},
    {`CALIPTRA_OWNER_PK_HASH_6_MASK,            `CALIPTRA_OWNER_PK_HASH_6,            `CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_6},
    {`CALIPTRA_OWNER_PK_HASH_7_MASK,            `CALIPTRA_OWNER_PK_HASH_7,            `CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_7},
    {`CALIPTRA_OWNER_PK_HASH_8_MASK,            `CALIPTRA_OWNER_PK_HASH_8,            `CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_8},
    {`CALIPTRA_OWNER_PK_HASH_9_MASK,            `CALIPTRA_OWNER_PK_HASH_9,            `CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_9},
    {`CALIPTRA_OWNER_PK_HASH_10_MASK,           `CALIPTRA_OWNER_PK_HASH_10,           `CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_10},
    {`CALIPTRA_OWNER_PK_HASH_11_MASK,           `CALIPTRA_OWNER_PK_HASH_11,           `CLP_SOC_IFC_REG_FUSE_OWNER_PK_HASH_11},
    {`CALIPTRA_KEY_MANIFEST_SVN_MASK,           `CALIPTRA_KEY_MANIFEST_SVN,           `CLP_SOC_IFC_REG_FUSE_FMC_KEY_MANIFEST_SVN},
    {`CALIPTRA_RUNTIME_SVN_0_MASK,              `CALIPTRA_RUNTIME_SVN_0,              `CLP_SOC_IFC_REG_FUSE_RUNTIME_SVN_0},
    {`CALIPTRA_RUNTIME_SVN_1_MASK,              `CALIPTRA_RUNTIME_SVN_1,              `CLP_SOC_IFC_REG_FUSE_RUNTIME_SVN_1},
    {`CALIPTRA_RUNTIME_SVN_2_MASK,              `CALIPTRA_RUNTIME_SVN_2,              `CLP_SOC_IFC_REG_FUSE_RUNTIME_SVN_2},
    {`CALIPTRA_RUNTIME_SVN_3_MASK,              `CALIPTRA_RUNTIME_SVN_3,              `CLP_SOC_IFC_REG_FUSE_RUNTIME_SVN_3},
    {`CALIPTRA_PUBLIC_SERIAL_NUMBER_0_MASK,     `CALIPTRA_PUBLIC_SERIAL_NUMBER_0,     `CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_7},
    {`CALIPTRA_PUBLIC_SERIAL_NUMBER_1_MASK,     `CALIPTRA_PUBLIC_SERIAL_NUMBER_1,     `CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_8},
    {`CALIPTRA_PUBLIC_SERIAL_NUMBER_2_MASK,     `CALIPTRA_PUBLIC_SERIAL_NUMBER_2,     `CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_9},
    {`CALIPTRA_PUBLIC_SERIAL_NUMBER_3_MASK,     `CALIPTRA_PUBLIC_SERIAL_NUMBER_3,     `CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_10},
    {`CALIPTRA_LMS_KEY_REVOKE_MASK_MASK,        `CALIPTRA_LMS_KEY_REVOKE_MASK,        `CLP_SOC_IFC_REG_FUSE_LMS_REVOCATION},
    {`CALIPTRA_FPF_TRNG_0_MASK,                 `CALIPTRA_FPF_TRNG_0,                 `CLP_SOC_IFC_REG_CPTRA_ITRNG_ENTROPY_CONFIG_0},
    {`CALIPTRA_FPF_TRNG_1_MASK,                 `CALIPTRA_FPF_TRNG_1,                 `CLP_SOC_IFC_REG_CPTRA_ITRNG_ENTROPY_CONFIG_1},
    {`CALIPTRA_HW_ID_MASK,                      `CALIPTRA_HW_ID,                      `CLP_SOC_IFC_REG_FUSE_SOC_STEPPING_ID},
    {`CALIPTRA_ANTI_ROLLBACK_DISABLE_MASK,      `CALIPTRA_ANTI_ROLLBACK_DISABLE,      `CLP_SOC_IFC_REG_FUSE_ANTI_ROLLBACK_DISABLE},
    {`CALIPTRA_KEY_MANIFEST_PK_HASH_MASK_MASK,  `CALIPTRA_KEY_MANIFEST_PK_HASH_MASK,  `CLP_SOC_IFC_REG_FUSE_KEY_MANIFEST_PK_HASH_MASK},
    {`CALIPTRA_LMS_VERIFY_ENABLE_MASK,          `CALIPTRA_LMS_VERIFY_ENABLE,          `CLP_SOC_IFC_REG_FUSE_LMS_VERIFY},
    {`CALIPTRA_IDEVID_CSR_REQUEST_MASK,         `CALIPTRA_IDEVID_CSR_REQUEST,         `CLP_SOC_IFC_REG_CPTRA_DBG_MANUF_SERVICE_REG},
    {`CALIPTRA_CERT_ATTRIB_RATS_MASK,           `CALIPTRA_CERT_ATTRIB_RATS,           `CLP_SOC_IFC_REG_FUSE_IDEVID_CERT_ATTR_6},
    {`CALIPTRA_SET_FUSE_DONE_MASK,              `CALIPTRA_SET_FUSE_DONE,              `CLP_SOC_IFC_REG_CPTRA_FUSE_WR_DONE},
    {32'hFFFF_FFFF,                             32'hFFFF_FFFF,                        32'hFFFF_FFFF}  //EOF
  };
  
  reg [$bits(fuse_lut_element_t)-1:0] rdata0q;

  always_ff @(posedge i_clk) begin
    if (i_readen) begin
      rdata0q <= FUSE_LUT[i_raddr];
    end
  end

  assign o_rdata = rdata0q;
  

endmodule

